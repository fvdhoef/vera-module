`default_nettype none

module composer(
    input  wire        rst,
    input  wire        clk,

    // Register interface
    input  wire  [4:0] regs_addr,
    input  wire  [7:0] regs_wrdata,
    output reg   [7:0] regs_rddata,
    input  wire        regs_write,

    // Layer 1 interface
    output wire  [8:0] layer1_line_idx,
    output wire        layer1_line_render_start,
    input  wire        layer1_line_render_done,
    input  wire        layer1_enabled,
    output wire  [9:0] layer1_lb_rdidx,
    input  wire  [7:0] layer1_lb_rddata,

    // Layer 2 interface
    output wire  [8:0] layer2_line_idx,
    output wire        layer2_line_render_start,
    input  wire        layer2_line_render_done,
    input  wire        layer2_enabled,
    output wire  [9:0] layer2_lb_rdidx,
    input  wire  [7:0] layer2_lb_rddata,

    // Sprite interface
    output wire  [8:0] sprites_line_idx,
    output wire        sprites_line_render_start,
    input  wire        sprites_line_render_done,
    input  wire        sprites_enabled,
    output wire  [9:0] sprites_lb_rdidx,
    input  wire [15:0] sprites_lb_rddata,
    output reg   [9:0] sprites_lb_wridx,
    output wire [15:0] sprites_lb_wrdata,
    output reg         sprites_lb_wren,

    // Display interface
    input  wire        display_next_frame,
    input  wire        display_next_line,
    input  wire        display_next_pixel,
    input  wire        display_current_field,
    output reg   [7:0] display_data,
    
    // Video selection
    output wire  [1:0] display_mode,
    output wire        chroma_disable);

    // MODE:
    // 0 - disabled, no video
    // 1 - VGA
    // 2 - NTSC video
    // 3 - RGB interlaced, composite sync (via VGA connector)

    //////////////////////////////////////////////////////////////////////////
    // Register interface
    //////////////////////////////////////////////////////////////////////////

    // CTRL0
    reg  [1:0] reg_mode_r;
    reg        chroma_disable_r;
    reg  [7:0] frac_x_incr_r;
    reg  [7:0] frac_y_incr_r;

    // Register interface read data
    always @* begin
        case (regs_addr)
            5'h0: regs_rddata = {5'b0, chroma_disable_r, reg_mode_r};
            5'h1: regs_rddata = frac_x_incr_r;
            5'h2: regs_rddata = frac_y_incr_r;
            default: regs_rddata = 8'h00;
        endcase
    end

    // Register interface write data
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            reg_mode_r          <= 2'd0;
            chroma_disable_r    <= 0;
            frac_x_incr_r       <= 8'd128;
            frac_y_incr_r       <= 8'd128;

        end else begin
            if (regs_write) begin
                case (regs_addr[3:0])
                    5'h0: begin
                        reg_mode_r       <= regs_wrdata[1:0];
                        chroma_disable_r <= regs_wrdata[2];
                    end
                    5'h1: begin
                        frac_x_incr_r    <= regs_wrdata;
                    end
                    5'h2: begin
                        frac_y_incr_r    <= regs_wrdata;
                    end
                endcase
            end
        end
    end

    wire [7:0] frac_x_incr = reg_mode_r[1] ? {1'b0, frac_x_incr_r[7:1]} : frac_x_incr_r;

    assign display_mode = reg_mode_r;
    assign chroma_disable = chroma_disable_r;

    //////////////////////////////////////////////////////////////////////////
    // Composer
    //////////////////////////////////////////////////////////////////////////
    reg [16:0] x_counter_r;
    wire [9:0] x_counter = x_counter_r[16:7];

    reg [15:0] y_counter_r;
    wire [8:0] y_counter = y_counter_r[15:7];

    reg render_start_r;
    always @(posedge clk) render_start_r <= display_next_line;

    // Output control signals to other units
    assign layer1_line_idx           = y_counter;
    assign layer1_line_render_start  = render_start_r;
    assign layer2_line_idx           = y_counter;
    assign layer2_line_render_start  = render_start_r;
    assign sprites_line_idx          = y_counter;
    assign sprites_line_render_start = render_start_r;
    assign layer1_lb_rdidx           = x_counter;
    assign layer2_lb_rdidx           = x_counter;
    assign sprites_lb_rdidx          = x_counter;

    assign sprites_lb_wrdata = 16'h0000;

    wire layer1_opaque = layer1_lb_rddata[7:0] != 8'h0;
    wire layer2_opaque = layer2_lb_rddata[7:0] != 8'h0;
    wire sprite_opaque = sprites_lb_rddata[7:0] != 8'h0;

    wire sprite_z1 = sprites_lb_rddata[9:8] != 2'd1;
    wire sprite_z2 = sprites_lb_rddata[9:8] != 2'd2;
    wire sprite_z3 = sprites_lb_rddata[9:8] != 2'd3;

    always @* begin
        display_data = 8'h00;
        if (sprites_enabled && sprite_opaque && sprite_z1) display_data = sprites_lb_rddata[7:0];
        if (layer1_enabled  && layer1_opaque)              display_data = layer1_lb_rddata;
        if (sprites_enabled && sprite_opaque && sprite_z2) display_data = sprites_lb_rddata[7:0];
        if (layer2_enabled  && layer2_opaque)              display_data = layer2_lb_rddata;
        if (sprites_enabled && sprite_opaque && sprite_z3) display_data = sprites_lb_rddata[7:0];
    end

    // Vertical counter
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            y_counter_r <= 'd0;

        end else begin
            if (display_next_line && y_counter < 'd480) begin
                y_counter_r <= y_counter_r + (reg_mode_r[1] ? {7'b0, frac_y_incr_r, 1'b0} : {8'b0, frac_y_incr_r});
            end

            if (display_next_frame) begin
                y_counter_r <= (reg_mode_r[1] && !display_current_field) ? {8'b0, frac_y_incr_r} : 'd0;
            end
        end
    end

    // Horizontal counter
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            x_counter_r <= 'd0;

            sprites_lb_wren  <= 0;
            sprites_lb_wridx <= 0;

        end else begin
            sprites_lb_wren <= 0;

            if (display_next_pixel && x_counter < 'd640) begin
                x_counter_r <= x_counter_r + frac_x_incr;

                sprites_lb_wridx <= x_counter;
                sprites_lb_wren  <= 1;
            end
            
            if (display_next_line) begin
                x_counter_r <= 0;
            end
        end
    end

endmodule
