`default_nettype none

module logsin_table(
    input  wire        clk,
    input  wire  [7:0] addr,
    output reg  [11:0] value) /* synthesis syn_romstyle = "EBR" */;

    reg [7:0] addr_r;
    always @(posedge(clk)) addr_r <= addr;

    always @* case (addr_r)
        8'd0: value <= 12'd2137;
        8'd1: value <= 12'd1731;
        8'd2: value <= 12'd1543;
        8'd3: value <= 12'd1419;
        8'd4: value <= 12'd1326;
        8'd5: value <= 12'd1252;
        8'd6: value <= 12'd1190;
        8'd7: value <= 12'd1137;
        8'd8: value <= 12'd1091;
        8'd9: value <= 12'd1050;
        8'd10: value <= 12'd1013;
        8'd11: value <= 12'd979;
        8'd12: value <= 12'd949;
        8'd13: value <= 12'd920;
        8'd14: value <= 12'd894;
        8'd15: value <= 12'd869;
        8'd16: value <= 12'd846;
        8'd17: value <= 12'd825;
        8'd18: value <= 12'd804;
        8'd19: value <= 12'd785;
        8'd20: value <= 12'd767;
        8'd21: value <= 12'd749;
        8'd22: value <= 12'd732;
        8'd23: value <= 12'd717;
        8'd24: value <= 12'd701;
        8'd25: value <= 12'd687;
        8'd26: value <= 12'd672;
        8'd27: value <= 12'd659;
        8'd28: value <= 12'd646;
        8'd29: value <= 12'd633;
        8'd30: value <= 12'd621;
        8'd31: value <= 12'd609;
        8'd32: value <= 12'd598;
        8'd33: value <= 12'd587;
        8'd34: value <= 12'd576;
        8'd35: value <= 12'd566;
        8'd36: value <= 12'd556;
        8'd37: value <= 12'd546;
        8'd38: value <= 12'd536;
        8'd39: value <= 12'd527;
        8'd40: value <= 12'd518;
        8'd41: value <= 12'd509;
        8'd42: value <= 12'd501;
        8'd43: value <= 12'd492;
        8'd44: value <= 12'd484;
        8'd45: value <= 12'd476;
        8'd46: value <= 12'd468;
        8'd47: value <= 12'd461;
        8'd48: value <= 12'd453;
        8'd49: value <= 12'd446;
        8'd50: value <= 12'd439;
        8'd51: value <= 12'd432;
        8'd52: value <= 12'd425;
        8'd53: value <= 12'd418;
        8'd54: value <= 12'd411;
        8'd55: value <= 12'd405;
        8'd56: value <= 12'd399;
        8'd57: value <= 12'd392;
        8'd58: value <= 12'd386;
        8'd59: value <= 12'd380;
        8'd60: value <= 12'd375;
        8'd61: value <= 12'd369;
        8'd62: value <= 12'd363;
        8'd63: value <= 12'd358;
        8'd64: value <= 12'd352;
        8'd65: value <= 12'd347;
        8'd66: value <= 12'd341;
        8'd67: value <= 12'd336;
        8'd68: value <= 12'd331;
        8'd69: value <= 12'd326;
        8'd70: value <= 12'd321;
        8'd71: value <= 12'd316;
        8'd72: value <= 12'd311;
        8'd73: value <= 12'd307;
        8'd74: value <= 12'd302;
        8'd75: value <= 12'd297;
        8'd76: value <= 12'd293;
        8'd77: value <= 12'd289;
        8'd78: value <= 12'd284;
        8'd79: value <= 12'd280;
        8'd80: value <= 12'd276;
        8'd81: value <= 12'd271;
        8'd82: value <= 12'd267;
        8'd83: value <= 12'd263;
        8'd84: value <= 12'd259;
        8'd85: value <= 12'd255;
        8'd86: value <= 12'd251;
        8'd87: value <= 12'd248;
        8'd88: value <= 12'd244;
        8'd89: value <= 12'd240;
        8'd90: value <= 12'd236;
        8'd91: value <= 12'd233;
        8'd92: value <= 12'd229;
        8'd93: value <= 12'd226;
        8'd94: value <= 12'd222;
        8'd95: value <= 12'd219;
        8'd96: value <= 12'd215;
        8'd97: value <= 12'd212;
        8'd98: value <= 12'd209;
        8'd99: value <= 12'd205;
        8'd100: value <= 12'd202;
        8'd101: value <= 12'd199;
        8'd102: value <= 12'd196;
        8'd103: value <= 12'd193;
        8'd104: value <= 12'd190;
        8'd105: value <= 12'd187;
        8'd106: value <= 12'd184;
        8'd107: value <= 12'd181;
        8'd108: value <= 12'd178;
        8'd109: value <= 12'd175;
        8'd110: value <= 12'd172;
        8'd111: value <= 12'd169;
        8'd112: value <= 12'd167;
        8'd113: value <= 12'd164;
        8'd114: value <= 12'd161;
        8'd115: value <= 12'd159;
        8'd116: value <= 12'd156;
        8'd117: value <= 12'd153;
        8'd118: value <= 12'd151;
        8'd119: value <= 12'd148;
        8'd120: value <= 12'd146;
        8'd121: value <= 12'd143;
        8'd122: value <= 12'd141;
        8'd123: value <= 12'd138;
        8'd124: value <= 12'd136;
        8'd125: value <= 12'd134;
        8'd126: value <= 12'd131;
        8'd127: value <= 12'd129;
        8'd128: value <= 12'd127;
        8'd129: value <= 12'd125;
        8'd130: value <= 12'd122;
        8'd131: value <= 12'd120;
        8'd132: value <= 12'd118;
        8'd133: value <= 12'd116;
        8'd134: value <= 12'd114;
        8'd135: value <= 12'd112;
        8'd136: value <= 12'd110;
        8'd137: value <= 12'd108;
        8'd138: value <= 12'd106;
        8'd139: value <= 12'd104;
        8'd140: value <= 12'd102;
        8'd141: value <= 12'd100;
        8'd142: value <= 12'd98;
        8'd143: value <= 12'd96;
        8'd144: value <= 12'd94;
        8'd145: value <= 12'd92;
        8'd146: value <= 12'd91;
        8'd147: value <= 12'd89;
        8'd148: value <= 12'd87;
        8'd149: value <= 12'd85;
        8'd150: value <= 12'd83;
        8'd151: value <= 12'd82;
        8'd152: value <= 12'd80;
        8'd153: value <= 12'd78;
        8'd154: value <= 12'd77;
        8'd155: value <= 12'd75;
        8'd156: value <= 12'd74;
        8'd157: value <= 12'd72;
        8'd158: value <= 12'd70;
        8'd159: value <= 12'd69;
        8'd160: value <= 12'd67;
        8'd161: value <= 12'd66;
        8'd162: value <= 12'd64;
        8'd163: value <= 12'd63;
        8'd164: value <= 12'd62;
        8'd165: value <= 12'd60;
        8'd166: value <= 12'd59;
        8'd167: value <= 12'd57;
        8'd168: value <= 12'd56;
        8'd169: value <= 12'd55;
        8'd170: value <= 12'd53;
        8'd171: value <= 12'd52;
        8'd172: value <= 12'd51;
        8'd173: value <= 12'd49;
        8'd174: value <= 12'd48;
        8'd175: value <= 12'd47;
        8'd176: value <= 12'd46;
        8'd177: value <= 12'd45;
        8'd178: value <= 12'd43;
        8'd179: value <= 12'd42;
        8'd180: value <= 12'd41;
        8'd181: value <= 12'd40;
        8'd182: value <= 12'd39;
        8'd183: value <= 12'd38;
        8'd184: value <= 12'd37;
        8'd185: value <= 12'd36;
        8'd186: value <= 12'd35;
        8'd187: value <= 12'd34;
        8'd188: value <= 12'd33;
        8'd189: value <= 12'd32;
        8'd190: value <= 12'd31;
        8'd191: value <= 12'd30;
        8'd192: value <= 12'd29;
        8'd193: value <= 12'd28;
        8'd194: value <= 12'd27;
        8'd195: value <= 12'd26;
        8'd196: value <= 12'd25;
        8'd197: value <= 12'd24;
        8'd198: value <= 12'd23;
        8'd199: value <= 12'd23;
        8'd200: value <= 12'd22;
        8'd201: value <= 12'd21;
        8'd202: value <= 12'd20;
        8'd203: value <= 12'd20;
        8'd204: value <= 12'd19;
        8'd205: value <= 12'd18;
        8'd206: value <= 12'd17;
        8'd207: value <= 12'd17;
        8'd208: value <= 12'd16;
        8'd209: value <= 12'd15;
        8'd210: value <= 12'd15;
        8'd211: value <= 12'd14;
        8'd212: value <= 12'd13;
        8'd213: value <= 12'd13;
        8'd214: value <= 12'd12;
        8'd215: value <= 12'd12;
        8'd216: value <= 12'd11;
        8'd217: value <= 12'd10;
        8'd218: value <= 12'd10;
        8'd219: value <= 12'd9;
        8'd220: value <= 12'd9;
        8'd221: value <= 12'd8;
        8'd222: value <= 12'd8;
        8'd223: value <= 12'd7;
        8'd224: value <= 12'd7;
        8'd225: value <= 12'd7;
        8'd226: value <= 12'd6;
        8'd227: value <= 12'd6;
        8'd228: value <= 12'd5;
        8'd229: value <= 12'd5;
        8'd230: value <= 12'd5;
        8'd231: value <= 12'd4;
        8'd232: value <= 12'd4;
        8'd233: value <= 12'd4;
        8'd234: value <= 12'd3;
        8'd235: value <= 12'd3;
        8'd236: value <= 12'd3;
        8'd237: value <= 12'd2;
        8'd238: value <= 12'd2;
        8'd239: value <= 12'd2;
        8'd240: value <= 12'd2;
        8'd241: value <= 12'd1;
        8'd242: value <= 12'd1;
        8'd243: value <= 12'd1;
        8'd244: value <= 12'd1;
        8'd245: value <= 12'd1;
        8'd246: value <= 12'd1;
        8'd247: value <= 12'd1;
        8'd248: value <= 12'd0;
        8'd249: value <= 12'd0;
        8'd250: value <= 12'd0;
        8'd251: value <= 12'd0;
        8'd252: value <= 12'd0;
        8'd253: value <= 12'd0;
        8'd254: value <= 12'd0;
        8'd255: value <= 12'd0;
    endcase

endmodule
